--
-- Author : Team G4

-- Design Unit: test_bench for 8x8 array multiplier, with verifier.


-- Revision History
-- Version 1.0
-- Date: 01-12-2022

--****************************************************
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity tb_array_8x8_mult is
end tb_array_8x8_mult;


architecture tb_array_8x8_mult_arch of tb_array_8x8_mult is

type test_vector_8x8_mult is record
  
  a: std_logic_vector(7 downto 0);
  b: std_logic_vector(7 downto 0);
  res: std_logic_vector(15 downto 0);
end record;

type test_vector_data is array (natural range <>) of test_vector_8x8_mult;

constant data_array: test_vector_data(57 downto 0) := 
(("00000010","00000001","0000000000000010"),
("00000010","00000010","0000000000000100"),
("11111111","10110011","1011001001001101"),
("10101010","11110000","1001111101100000"),
("00000010","00000101","0000000000001010"),
("00000010","00000110","0000000000001100"),
("00000010","00000111","0000000000001110"),
("00000010","00001000","0000000000010000"),
("00000010","00001001","0000000000010010"),
("00000010","00001010","0000000000010100"),
("00000010","00001011","0000000000010110"),
("00000010","00001100","0000000000011000"),
("00000010","00001101","0000000000011010"),
("00000010","00001110","0000000000011100"),
("00000010","00001111","0000000000011110"),
("00010110","01000101","0000010111101110"),
("01000101","00101010","0000101101010010"),
("01100000","00111001","0001010101100000"),
("01100001","01010100","0001111111010100"),
("00000100","00010100","0000000001010000"),
("01011001","00001001","0000001100100001"),
("01000010","00100111","0000101000001110"),
("00010110","01000010","0000010110101100"),
("00111010","00000010","0000000001110100"),
("00110110","01011111","0001010000001010"),
("01000010","01001101","0001001111011010"),
("01000111","01010001","0001011001110111"),
("00000110","00001010","0000000000111100"),
("00110111","01000000","0000110111000000"),
("00111110","01011000","0001010101010000"),
("01100011","01000110","0001101100010010"),
("00011001","00011010","0000001010001010"),
("01010010","00110100","0001000010101000"),
("00111011","00110101","0000110000110111"),
("01011001","00001110","0000010011011110"),
("00011101","01011101","0000101010001001"),
("01110011","11011110","0110001110111010"),
("01110100","11101010","0110101000001000"),
("01110101","11100010","0110011101001010"),
("01110110","11101000","0110101011110000"),
("01110111","10011100","0100100010000100"),
("01111000","11101001","0110110100111000"),
("10100101","11110100","1001110101000100"),
("10101000","11111001","1010001101101000"),
("10101001","11111100","1010011001011100"),
("10100010","11111010","1001111000110100"),
("10100110","11011100","1000111010101000"),
("10101011","10110001","0111011000111011"),
("10101110","10110100","0111101001011000"),
("10100100","10100000","0110011010000000"),
("10110010","11111110","1011000010011100"),
("10101111","10100011","0110111101101101"),
("01111100","10111110","0101110000001000"),
("01111111","11000100","0110000100111100"),
("01111011","11111011","0111100010011001"),
("01111101","11100111","0111000011001011"),
("10000001","11101101","0111011101101101"),
("11111111","11111111","1111111000000001"));

component array_multiplier_8bit is
  Port ( 
  A : in std_logic_vector (7 downto 0);
  B : in std_logic_vector (7 downto 0);
  Z : out std_logic_vector (15 downto 0));
end component;

signal a_test, b_test: std_logic_vector(7 downto 0);
signal res_test: std_logic_vector(15 downto 0);
signal test_ok: boolean;

begin
  uut:array_multiplier_8bit
  port map(A=>a_test, B=>b_test, Z=>res_test);
    
    process begin
      for i in data_array'range loop
        a_test <= data_array(i).a;
        b_test <= data_array(i).b;
        wait for 10 ns;
        if res_test /= data_array(i).res then
          test_ok <= FALSE;
        else
          test_ok <= TRUE;
        end if;
      end loop;
      wait;
    end process;
  end tb_array_8x8_mult_arch;
