library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity tb_expression_calculator_top_level is
end tb_expression_calculator_top_level;


architecture tb_expression_calculator_top_level_arch of tb_expression_calculator_top_level is

type test_vector_toplevel is record
  
  a: std_logic_vector(7 downto 0);
  b: std_logic_vector(7 downto 0);
  res: signed(15 downto 0);
  load_in : std_logic;
  load_out :std_logic;
end record;

type test_vector_data is array (natural range <>) of test_vector_toplevel;

constant data_array: test_vector_data(67 downto 0) := 
(("00001000","00000101","0000000000001011",'1','1'),
("00000010","00001010","0000000000000110",'1','1'),
("10101010","11001100","0010000111011111",'1','1'),
("00011101","01011101","0010000111011111",'0','0'),    -- when input Load is 0, inputs are changed but output remains the same as previous
("00001111","00010110","0000000001010011",'1','1'),
("00010000","00100010","0000000010001001",'1','1'),
("00010001","00011010","0000000001101111",'1','1'),
("00010010","00100000","0000000010010001",'1','1'),
("00010011","00111000","0000000100001011",'1','1'),
("00010100","00100001","0000000010100110",'1','1'),
("01000001","00101100","0000001011001100",'1','1'),
("01000100","00110001","0000001101000010",'1','1'),
("01000101","00110100","0000001110000010",'1','1'),
("00111110","00110010","0000001100001000",'1','1'),
("01000010","00010100","0000000101001011",'1','1'),
("01000111","01001101","0000010101010111",'1','1'),
("01001010","01010000","0000010111001001",'1','1'),
("01000000","00111100","0000001111000001",'1','1'),
("01001110","00110110","0000010000011110",'1','1'),
("01001011","00111111","0000010010011110",'1','1'),
("00011000","01011010","0000001000011101",'1','1'),
("00011011","01100000","0000001010001001",'1','1'),
("00010111","01100100","0000001001000000",'1','1'),
("00011001","01100011","0000001001101011",'1','1'),
("00011101","01011101","0000001010100011",'1','1'),
("00010110","01000101","0000000101111100",'1','1'),
("01000101","00101010","0000001011010101",'1','1'),
("01100000","00111001","0000010101011001",'1','1'),
("01100001","01010100","0000011111110110",'1','1'),
("00000100","00010100","0000000000010101",'1','1'),
("01011001","00001001","0000000011001001",'1','1'),
("01000010","00100111","0000001010000100",'1','1'),
("00010110","01000010","0000000101101100",'1','1'),
("00111010","00000010","0000000000011110",'1','1'),
("00110110","01011111","0000010100000011",'1','1'),
("01000010","01001101","0000010011110111",'1','1'),
("01000111","01010001","0000010110011110",'1','1'),
("00000110","00001010","0000000000010000",'1','1'),
("00110111","01000000","0000001101110001",'1','1'),
("00111110","01011000","0000010101010101",'1','1'),
("01100011","01000110","0000011011000101",'1','1'),
("00011001","00011010","0000011011000101",'1','1'),
("01010010","00110100","0000010000101011",'1','1'),
("00111011","00110101","0000001100001110",'1','1'),
("01011001","00001110","0000000100111000",'1','1'),
("00011101","01011101","0000001010100011",'1','1'),
("01110011","11011110","0001100011101111",'1','1'),
("01110100","11101010","0001101010000011",'1','1'),
("01110101","11100010","0001100111010011",'1','1'),
("01110110","11101000","0001101010111101",'1','1'),
("01110111","10011100","0001001000100010",'1','1'),
("01111000","11101001","0001101101001111",'1','1'),
("10100101","11110100","0010011101010010",'1','1'),
("10101000","11111001","0010100011011011",'1','1'),
("10101001","11111100","0010100110011000",'1','1'),
("10100010","11111010","0010011110001110",'1','1'),
("10100110","11011100","0010001110101011",'1','1'),
("10101011","10110001","0001110110001111",'1','1'),
("10101110","10110100","0001111010010111",'1','1'),
("10100100","10100000","0001100110100001",'1','1'),
("10110010","11111110","0010110000101000",'1','1'),
("10101111","10100011","0001101111011100",'1','1'),
("01111100","10111110","0001011100000011",'1','1'),
("01111111","11000100","0001100001010000",'1','1'),
("01111011","11111011","0001111000100111",'1','1'),
("01111101","11100111","0001110000110011",'1','1'),
("10000001","11101101","0001110111011100",'1','1'),
("11111111","11111111","0011111110000001",'1','1'));  

component expression_calculator_top_level is
  port(
    A, B: in std_logic_vector(7 downto 0);
    clk, rst, load_in, load_out: in std_logic;
    end_flag: out std_logic;
    Z: out signed(15 downto 0));
    
  end component;

signal a_test, b_test: std_logic_vector(7 downto 0) := (others=>'0');
signal res_test: signed(15 downto 0) := (others=>'0');
signal test_clk, test_rst, test_load_in,test_load_out, test_endflag: std_logic := '0';

signal test_ok: boolean;

begin
  
  --Clock pulses
  clock:process
  begin
    wait for 10 ns;
          test_clk <= '1';
          wait for 10 ns;
          test_clk <= '0';
    end process clock;
    
    
    
  uut:expression_calculator_top_level
  port map(A=>a_test, B=>b_test,clk=>test_clk,rst=>test_rst,load_in=>test_load_in,load_out=>test_load_out,end_flag=>test_endflag, Z=>res_test);
    
    process 
     begin
       
       -- Reset the system--
       test_rst <= '1';
      wait for 40 ns;
       test_rst <= '0';
      wait for 20 ns;
      
      for i in data_array'range loop
        test_load_in <= data_array(i).load_in;
        a_test <= data_array(i).a;
        b_test <= data_array(i).b;
        wait for 30 ns;
        test_load_out <= data_array(i).load_out;
        wait for 30 ns;
        if res_test /= data_array(i).res then
          test_ok <= FALSE;
        else
          test_ok <= TRUE;
        end if;
        test_load_out <= '0';
      end loop;
      wait;
    end process;
  end tb_expression_calculator_top_level_arch;
